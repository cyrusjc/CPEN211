module lab8_top(KEY,SW,LEDR,HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,CLOCK_50);
	
	`define MREAD 2'b00
	`define MWRITE 2'b01

	input [3:0] KEY;
	input [9:0] SW;
	output [9:0] LEDR;
	output [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
	input CLOCK_50;
	
	wire clk = CLOCK_50;
	wire reset = ~KEY[1];
	wire s = ~KEY[2];
	wire load = ~KEY[3];

	wire [15:0] x; //X IS AN INPUT FROM MEM (TO IREG)
	wire [1:0] mem_cmd;
	wire [8:0] mem_addr;
	wire [15:0] out; // OUT ALSO GOES TO MEM DIN
	//INSTANTIATING CPU
	cpu CPU(clk,reset,x,out,N,V,Z,mem_cmd,mem_addr,LEDR[8]);
	

	wire [15:0] dout;
	wire msel = 1'b0 == mem_addr[8:8];
	wire isMREAD = `MREAD == mem_cmd; // WIRING STUFF TO SEE EASILY
	wire e = msel & isMREAD; // e IS INPUT TO TRISTATE
	assign x = e ? dout : 16'bz;
	wire isMWRITE = `MWRITE == mem_cmd;
	wire write = isMWRITE & msel;
	//INSTANTIATING MEM
	RAM MEM(clk,mem_addr[7:0],mem_addr[7:0],write,out,dout);

	//LAb 7: STAGE 3
	//INPUT THING
	wire [15:0] SWin = {6'b0,SW[9:0]};
	//wire [15:0] SWout;
	wire e1 = (mem_cmd == `MREAD) & (mem_addr == 9'b101000000);
	assign x = e1 ? SWin : 16'bz;

	//OUTPUT
	//wire LEDRin [7:0] = out[7:0];
	wire e2 = (mem_cmd == `MWRITE) & (mem_addr == 9'b100000000);
	vDFFE #(8) ledREG(clk,e2,out[7:0],LEDR[7:0]);

	assign HEX0 = 7'b1111111;
	assign HEX1 = 7'b1111111;
	assign HEX2 = 7'b1111111;
	assign HEX3 = 7'b1111111;
	assign HEX4 = 7'b1111111;
	assign HEX5 = 7'b1111111;
	assign LEDR[9] = 1'b0;

	
endmodule


module RAM(clk,read_address,write_address,write,din,dout);
	parameter data_width = 16;
	parameter addr_width = 8;
	parameter filename = "lab8fig2.txt";
	
	input 		clk;
	input 		[addr_width-1:0] read_address, write_address;
	input 		write;
	input 		[data_width-1:0] din;
	output reg 	[data_width-1:0] dout;

	reg [data_width-1:0] mem [2**addr_width-1:0];

	initial $readmemb(filename,mem);

	always @(posedge clk) begin
		if(write)
			mem[write_address] <= din;
		dout <= mem[read_address];
	end
endmodule
